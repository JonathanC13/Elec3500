** Profile: "SCHEMATIC1-SimNMOS2"  [ P:\CourseNotes\ELEC3500\Lab1_2005\nmos2-schematic1-simnmos2.sim ] 

** Creating circuit file "nmos2-schematic1-simnmos2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\nmos2.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 120ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\nmos2-SCHEMATIC1.net" 


.END
