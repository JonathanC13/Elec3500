** Profile: "SCHEMATIC1-SimNMOS1"  [ W:\ELEC3500\lab1\Lab1_2006\1\nmos1-pspicefiles\schematic1\simnmos1.sim ] 

** Creating circuit file "SimNMOS1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../nmos1-pspicefiles/nmos1.lib" 
* From [PSPICE NETLIST] section of W:\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 0 5 0.5 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
