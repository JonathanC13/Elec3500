** Profile: "SCHEMATIC1-SimNMOS1"  [ P:\CourseNotes\ELEC3500\Lab1_2005\nmos1-schematic1-simnmos1.sim ] 

** Creating circuit file "nmos1-schematic1-simnmos1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\nmos1.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 120ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\nmos1-SCHEMATIC1.net" 


.END
