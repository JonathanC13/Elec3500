** Profile: "SCHEMATIC1-SimPMOS!"  [ P:\CourseNotes\ELEC3500\Lab1_2005\pmos1-schematic1-simpmos!.sim ] 

** Creating circuit file "pmos1-schematic1-simpmos!.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\pmos1.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 120ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pmos1-SCHEMATIC1.net" 


.END
